library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity valida_prod is
    port (
        
        
    );
end entity valida_prod;

architecture rtl of valida_prod is
    
begin
    
    
end architecture rtl;